
// Copyright (c) 2016 Massachusetts Institute of Technology

// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

/**
 * This package provides a collection of modules and interfaces for creating
 * and accessing SRAM cells. For FPGA and simulation targets, this package
 * uses the standard BRAM and BRAM_CORE packages. For ASIC targets, this
 * package can be used as placeholders for SRAMs generated by memory
 * compilers.
 */
package SRAMUtil;

import BRAMCore::*;
import RevertingVirtualReg::*;

import Ehr::*;

// If SRAMUTIL_SRAM is defined, then this package will use SRAM
//`define SRAMUTIL_SRAM

`ifdef SRAMUTIL_SRAM
import SRAMCore::*;
`endif

/// Single port SRAM interface
interface SRAM_1RW#(type addrT, type dataT);
    method Action req(Bool write, addrT a, dataT d);
    method dataT readData;
    method Action readDataDeq;
endinterface

/// Simple dual port SRAM interface (1 read port and 1 write port)
interface SRAM_1R1W#(type addrT, type dataT);
    // write port
    method Action writeReq(addrT a, dataT d);
    // read port
    method Action readReq(addrT a);
    method dataT readData;
    method Action readDataDeq;
endinterface

/// True dual port SRAM interface (2 read/write ports)
interface SRAM_2RW#(type addrT, type dataT);
    // port A
    interface SRAM_1RW#(addrT, dataT) a;
    // port B
    interface SRAM_1RW#(addrT, dataT) b;
endinterface

/**
 * Single-Port SRAM
 *
 * readData < readDataDeq < req
 */
module mkSRAM_1RW( SRAM_1RW#(addrT, dataT) ) provisos (Bits#(addrT, addrSz), Bits#(dataT, dataSz));
    Integer memSz = valueOf(TExp#(addrSz));
    Bool hasOutputRegister = False;
`ifdef SRAMUTIL_SRAM
    SRAMCore1RW#(addrT, dataT) sram <- mkSRAMCore1RW;
`else
    BRAM_PORT#(addrT, dataT) bram <- mkBRAMCore1(memSz, hasOutputRegister);
`endif

    Ehr#(2, Bool) readPending <- mkEhr(False);

    method Action req(Bool write, addrT a, dataT d) if (!readPending[1]);
`ifdef SRAMUTIL_SRAM
        sram.req(write, a, d);
`else
        bram.put(write, a, d);
`endif
        if (!write) begin
            readPending[1] <= True;
        end
    endmethod
    method dataT readData if (readPending[0]);
`ifdef SRAMUTIL_SRAM
        return sram.readData;
`else
        return bram.read;
`endif
    endmethod
    method Action readDataDeq;
        readPending[0] <= False;
    endmethod
endmodule

`ifdef SRAMUTIL_SRAM
module mkSRAM_1RW_64x52( SRAM_1RW#(Bit#(6), Bit#(52)) );
    Integer memSz = valueOf(TExp#(6));
    Bool hasOutputRegister = False;

    SRAMCore1RW#(Bit#(6), Bit#(52)) sram <- mkSRAMCore1RW_64x52;
    Ehr#(2, Bool) readPending <- mkEhr(False);

    method Action req(Bool write, Bit#(6) a, Bit#(52) d) if (!readPending[1]);
        sram.req(write, a, d);
        if (!write) begin
            readPending[1] <= True;
        end
    endmethod
    method Bit#(52) readData if (readPending[0]);
        return sram.readData;
    endmethod
    method Action readDataDeq;
        readPending[0] <= False;
    endmethod
endmodule

module mkSRAM_1RW_64x64( SRAM_1RW#(Bit#(6), Bit#(64)) );
    Integer memSz = valueOf(TExp#(6));
    Bool hasOutputRegister = False;

    SRAMCore1RW#(Bit#(6), Bit#(64)) sram <- mkSRAMCore1RW_64x64;
    Ehr#(2, Bool) readPending <- mkEhr(False);

    method Action req(Bool write, Bit#(6) a, Bit#(64) d) if (!readPending[1]);
        sram.req(write, a, d);
        if (!write) begin
            readPending[1] <= True;
        end
    endmethod
    method Bit#(64) readData if (readPending[0]);
        return sram.readData;
    endmethod
    method Action readDataDeq;
        readPending[0] <= False;
    endmethod
endmodule
`endif
/**
 * Simple Dual-Port SRAM
 *
 * A concurrent read and write to the same address will result in the read
 * seeing the *old* data.
 *
 * readData < readDataDeq < readReq < writeReq 
 */
module mkSRAM_1R1W( SRAM_1R1W#(addrT, dataT) ) provisos (Bits#(addrT, addrSz), Bits#(dataT, dataSz));
    Integer memSz = valueOf(TExp#(addrSz));
    Bool hasOutputRegister = False;
`ifdef SRAMUTIL_SRAM
    SRAMCore1R1W#(addrT, dataT) sram <- mkSRAMCore1R1W;
`else
    BRAM_DUAL_PORT#(addrT, dataT) bram <- mkBRAMCore2(memSz, hasOutputRegister);
`endif

    Ehr#(2, Bool) readPending <- mkEhr(False);
    Reg#(Bool) _rvr_readReq_sb_writeReq <- mkRevertingVirtualReg(True);

    method Action writeReq(addrT a, dataT d);
`ifdef SRAMUTIL_SRAM
        sram.writeReq(a, d);
`else
        bram.a.put(True, a, d);
`endif

        // reverting virtual register for scheduling purposes
        _rvr_readReq_sb_writeReq <= False;
    endmethod

    method Action readReq(addrT a) if (!readPending[1] && _rvr_readReq_sb_writeReq);
`ifdef SRAMUTIL_SRAM
        sram.readReq(a);
`else
        bram.b.put(False, a, unpack(0));
`endif
        readPending[1] <= True;
    endmethod
    method dataT readData if (readPending[0]);
`ifdef SRAMUTIL_SRAM
        return sram.readData;
`else
        return bram.b.read;
`endif
    endmethod
    method Action readDataDeq;
        readPending[0] <= False;
    endmethod
endmodule


/*module mkSRAM_1R1W_64x64( SRAM_1R1W#(addrT, dataT) ) provisos (Bits#(addrT, 6), Bits#(dataT, 64));
    Integer memSz = valueOf(TExp#(6));
    Bool hasOutputRegister = False;

    SRAMCore1R1W#(addrT, dataT) sram <- mkSRAMCore1R1W_64x64;

    Ehr#(2, Bool) readPending <- mkEhr(False);
    Reg#(Bool) _rvr_readReq_sb_writeReq <- mkRevertingVirtualReg(True);

    method Action writeReq(addrT a, dataT d);
        sram.writeReq(a, d);
        // reverting virtual register for scheduling purposes
        _rvr_readReq_sb_writeReq <= False;
    endmethod

    method Action readReq(addrT a) if (!readPending[1] && _rvr_readReq_sb_writeReq);

        sram.readReq(a);

        readPending[1] <= True;
    endmethod
    method dataT readData if (readPending[0]);
        return sram.readData;

    endmethod
    method Action readDataDeq;
        readPending[0] <= False;
    endmethod
endmodule


module mkSRAM_1R1W_64x52( SRAM_1R1W#(addrT, dataT) ) provisos (Bits#(addrT, 6), Bits#(dataT, 52));
    Integer memSz = valueOf(TExp#(6));
    Bool hasOutputRegister = False;

    SRAMCore1R1W#(addrT, dataT) sram <- mkSRAMCore1R1W_64x52;

    Ehr#(2, Bool) readPending <- mkEhr(False);
    Reg#(Bool) _rvr_readReq_sb_writeReq <- mkRevertingVirtualReg(True);

    method Action writeReq(addrT a, dataT d);
        sram.writeReq(a, d);
        // reverting virtual register for scheduling purposes
        _rvr_readReq_sb_writeReq <= False;
    endmethod

    method Action readReq(addrT a) if (!readPending[1] && _rvr_readReq_sb_writeReq);

        sram.readReq(a);

        readPending[1] <= True;
    endmethod
    method dataT readData if (readPending[0]);
        return sram.readData;

    endmethod
    method Action readDataDeq;
        readPending[0] <= False;
    endmethod
endmodule


module mkSRAM_1R1W_64x4( SRAM_1R1W#(addrT, dataT) ) provisos (Bits#(addrT, 6), Bits#(dataT, 2));
    Integer memSz = valueOf(TExp#(6));
    Bool hasOutputRegister = False;

    SRAMCore1R1W#(addrT, dataT) sram <- mkSRAMCore1R1W_64x2;

    Ehr#(2, Bool) readPending <- mkEhr(False);
    Reg#(Bool) _rvr_readReq_sb_writeReq <- mkRevertingVirtualReg(True);

    method Action writeReq(addrT a, dataT d);
        sram.writeReq(a, d);
        // reverting virtual register for scheduling purposes
        _rvr_readReq_sb_writeReq <= False;
    endmethod

    method Action readReq(addrT a) if (!readPending[1] && _rvr_readReq_sb_writeReq);

        sram.readReq(a);

        readPending[1] <= True;
    endmethod
    method dataT readData if (readPending[0]);
        return sram.readData;

    endmethod
    method Action readDataDeq;
        readPending[0] <= False;
    endmethod
endmodule*/

/**
 * Simple Dual-Port SRAM with bypassing
 *
 * A concurrent read and write to the same address will result in the read
 * seeing the *new* data.
 *
 * readData < readDataDeq < readReq
 * writeReq < readReq
 * writeReq CF {readData, readDataDeq}
 */
module mkSRAM_1R1W_Bypass( SRAM_1R1W#(addrT, dataT) ) provisos (Bits#(addrT, addrSz), Bits#(dataT, dataSz));
    Integer memSz = valueOf(TExp#(addrSz));
    Bool hasOutputRegister = False;
`ifdef SRAMUTIL_SRAM
    SRAMCore1R1W#(addrT, dataT) sram <- mkSRAMCore1R1W;
`else
    BRAM_DUAL_PORT#(addrT, dataT) bram <- mkBRAMCore2(memSz, hasOutputRegister);
`endif

    Ehr#(2, Bool) readPending <- mkEhr(False);
    Ehr#(2, Maybe#(dataT)) bypassData <- mkEhr(tagged Invalid);

    Wire#(Maybe#(Tuple2#(addrT, dataT))) writeReqWire <- mkDWire(tagged Invalid);

    method Action writeReq(addrT a, dataT d);
`ifdef SRAMUTIL_SRAM
        sram.writeReq(a, d);
`else
        bram.a.put(True, a, d);
`endif
        writeReqWire <= tagged Valid tuple2(a, d);
    endmethod

    method Action readReq(addrT a) if (!readPending[1]);
`ifdef SRAMUTIL_SRAM
        sram.readReq(a);
`else
        bram.b.put(False, a, unpack(0));
`endif
        readPending[1] <= True;
        if (writeReqWire matches tagged Valid {.writeAddr, .writeData} &&& pack(writeAddr) == pack(a)) begin
            bypassData[1] <= tagged Valid writeData;
        end
    endmethod
    method dataT readData if (readPending[0]);
        if (bypassData[0] matches tagged Valid .bypassData) begin
            return bypassData;
        end else begin
`ifdef SRAMUTIL_SRAM
            return sram.readData;
`else
            return bram.b.read;
`endif
        end
    endmethod
    method Action readDataDeq;
        readPending[0] <= False;
        if (isValid(bypassData[0])) begin
            bypassData[0] <= tagged Invalid;
        end
    endmethod
endmodule

`ifdef SRAMUTIL_SRAM
module mkSRAM_1R1W_Bypass_64x64( SRAM_1R1W#(Bit#(6), Bit#(64)) );
    Integer memSz = valueOf(TExp#(6));
    Bool hasOutputRegister = False;

    SRAMCore1R1W#(Bit#(6), Bit#(64)) sram <- mkSRAMCore1R1W_64x64;


    Ehr#(2, Bool) readPending <- mkEhr(False);
    Ehr#(2, Maybe#(Bit#(64))) bypassData <- mkEhr(tagged Invalid);

    Wire#(Maybe#(Tuple2#(Bit#(6), Bit#(64)))) writeReqWire <- mkDWire(tagged Invalid);

    method Action writeReq(Bit#(6) a, Bit#(64) d);

        sram.writeReq(a, d);

        writeReqWire <= tagged Valid tuple2(a, d);
    endmethod

    method Action readReq(Bit#(6) a) if (!readPending[1]);

        sram.readReq(a);

        readPending[1] <= True;
        if (writeReqWire matches tagged Valid {.writeAddr, .writeData} &&& pack(writeAddr) == pack(a)) begin
            bypassData[1] <= tagged Valid writeData;
        end
    endmethod
    method Bit#(64) readData if (readPending[0]);
        if (bypassData[0] matches tagged Valid .bypassData) begin
            return bypassData;
        end else begin
            return sram.readData;
        end
    endmethod
    method Action readDataDeq;
        readPending[0] <= False;
        if (isValid(bypassData[0])) begin
            bypassData[0] <= tagged Invalid;
        end
    endmethod
endmodule

module mkSRAM_1R1W_Bypass_64x52( SRAM_1R1W#(Bit#(6), Bit#(52)) );
    Integer memSz = valueOf(TExp#(6));
    Bool hasOutputRegister = False;

    SRAMCore1R1W#(Bit#(6), Bit#(52)) sram <- mkSRAMCore1R1W_64x52;


    Ehr#(2, Bool) readPending <- mkEhr(False);
    Ehr#(2, Maybe#(Bit#(52))) bypassData <- mkEhr(tagged Invalid);

    Wire#(Maybe#(Tuple2#(Bit#(6), Bit#(52)))) writeReqWire <- mkDWire(tagged Invalid);

    method Action writeReq(Bit#(6) a, Bit#(52) d);

        sram.writeReq(a, d);

        writeReqWire <= tagged Valid tuple2(a, d);
    endmethod

    method Action readReq(Bit#(6) a) if (!readPending[1]);

        sram.readReq(a);

        readPending[1] <= True;
        if (writeReqWire matches tagged Valid {.writeAddr, .writeData} &&& pack(writeAddr) == pack(a)) begin
            bypassData[1] <= tagged Valid writeData;
        end
    endmethod
    method Bit#(52) readData if (readPending[0]);
        if (bypassData[0] matches tagged Valid .bypassData) begin
            return bypassData;
        end else begin
            return sram.readData;
        end
    endmethod
    method Action readDataDeq;
        readPending[0] <= False;
        if (isValid(bypassData[0])) begin
            bypassData[0] <= tagged Invalid;
        end
    endmethod
endmodule

module mkSRAM_1R1W_Bypass_64x2( SRAM_1R1W#(Bit#(6), dataT) ) provisos (Bits#(dataT, 2));
    Integer memSz = valueOf(TExp#(6));
    Bool hasOutputRegister = False;

    SRAMCore1R1W#(Bit#(6), dataT) sram <- mkSRAMCore1R1W_64x2;


    Ehr#(2, Bool) readPending <- mkEhr(False);
    Ehr#(2, Maybe#(dataT)) bypassData <- mkEhr(tagged Invalid);

    Wire#(Maybe#(Tuple2#(Bit#(6), dataT))) writeReqWire <- mkDWire(tagged Invalid);

    method Action writeReq(Bit#(6) a, dataT d);

        sram.writeReq(a, d);

        writeReqWire <= tagged Valid tuple2(a, d);
    endmethod

    method Action readReq(Bit#(6) a) if (!readPending[1]);

        sram.readReq(a);

        readPending[1] <= True;
        if (writeReqWire matches tagged Valid {.writeAddr, .writeData} &&& pack(writeAddr) == pack(a)) begin
            bypassData[1] <= tagged Valid writeData;
        end
    endmethod
    method dataT readData if (readPending[0]);
        if (bypassData[0] matches tagged Valid .bypassData) begin
            return bypassData;
        end else begin
            return sram.readData;
        end
    endmethod
    method Action readDataDeq;
        readPending[0] <= False;
        if (isValid(bypassData[0])) begin
            bypassData[0] <= tagged Invalid;
        end
    endmethod
endmodule
`endif

/**
 * True Dual-Port SRAM.
 *
 * Has the additional constraint that a.req < b.req so that writes to port A
 * can be bypassed to reads from port B.
 */
module mkSRAM_2RW( SRAM_2RW#(addrT, dataT) ) provisos (Bits#(addrT, addrSz), Bits#(dataT, dataSz));
    Integer memSz = 0;
    Bool hasOutputRegister = False;
    BRAM_DUAL_PORT#(addrT, dataT) bram <- mkBRAMCore2(memSz, hasOutputRegister);

    Ehr#(2, Bool) readPendingA <- mkEhr(False);
    Ehr#(2, Bool) readPendingB <- mkEhr(False);

    // This is for bypassing writes to port A to reads from port B
    Ehr#(2, Maybe#(dataT)) bypassData <- mkEhr(tagged Invalid);
    Wire#(Maybe#(Tuple2#(addrT, dataT))) writeReqWire <- mkDWire(tagged Invalid);

    interface SRAM_1RW a;
        method Action req(Bool write, addrT a, dataT d) if (!readPendingA[1]);
            bram.a.put(write, a, d);
            if (!write) begin
                readPendingA[1] <= True;
            end else begin
                writeReqWire <= tagged Valid tuple2(a, d);
            end
        endmethod
        method dataT readData if (readPendingA[0]);
            return bram.a.read;
        endmethod
        method Action readDataDeq;
            readPendingA[0] <= False;
        endmethod
    endinterface
    interface SRAM_1RW b;
        method Action req(Bool write, addrT a, dataT d) if (!readPendingB[1]);
            bram.b.put(write, a, d);
            if (!write) begin
                readPendingB[1] <= True;
                if (writeReqWire matches tagged Valid {.writeAddr, .writeData} &&& pack(writeAddr) == pack(a)) begin
                    // bypassing from port A
                    bypassData[1] <= tagged Valid writeData;
                end
            end
        endmethod
        method dataT readData if (readPendingB[0]);
            if (bypassData[1] matches tagged Valid .bypass) begin
                return bypass;
            end else begin
                return bram.b.read;
            end
        endmethod
        method Action readDataDeq;
            readPendingB[0] <= False;
            if (isValid(bypassData[0])) begin
                bypassData[0] <= tagged Invalid;
            end
        endmethod
    endinterface
endmodule

endpackage
