// generated by gen_VerilogEHR.py using VerilogEHRWrapper.mako

// Copyright (c) 2019 Massachusetts Institute of Technology
//
// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

import Vector::*;

// This package uses Arrays for EHR interfaces in order to avoid needing
// a typeclass to say if there is an implementation of a VerilogEHR with
// the given number of ports.
typedef Array#(Reg#(t)) VerilogEHR#(type t);

(* always_ready *)
interface VerilogEHR_1_Raw#(numeric type dataSz);
    method Bit#(dataSz) read_0;
    method Action write_0(Bit#(dataSz) x);
endinterface

import "BVI" EHR_1 =
module mkVerilogEHR_1_Raw#(Bit#(dataSz) init)(VerilogEHR_1_Raw#(dataSz));
    parameter DATA_SZ = valueOf(dataSz);
    parameter RESET_VAL = init;

    default_clock clk(CLK);
    default_reset rst(RST_N);

    method read_0 read_0;
    method write_0(write_0) enable (EN_write_0);

    // intra-port scheduling
    schedule (read_0) CF (read_0);
    schedule (read_0) SB (write_0);
    schedule (write_0) SBR (write_0);

    // inter-port scheduling

    // paths
endmodule

import "BVI" EHRU_1 =
module mkVerilogEHRU_1_Raw(VerilogEHR_1_Raw#(dataSz));
    parameter DATA_SZ = valueOf(dataSz);

    default_clock clk(CLK);
    no_reset;

    method read_0 read_0;
    method write_0(write_0) enable (EN_write_0);

    // intra-port scheduling
    schedule (read_0) CF (read_0);
    schedule (read_0) SB (write_0);
    schedule (write_0) SBR (write_0);

    // inter-port scheduling

    // paths
endmodule

module mkVerilogEHR_1#(dataT init)(VerilogEHR#(dataT)) provisos (Bits#(dataT, dataSz));
    VerilogEHR_1_Raw#(dataSz) ehr_raw <- mkVerilogEHR_1_Raw(pack(init));
    Reg#(dataT) ehr_ifc[1];
    
    ehr_ifc[0] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_0);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_0(pack(x));
            endmethod
        endinterface);

    return ehr_ifc;
endmodule

module mkVerilogEHRU_1(VerilogEHR#(dataT)) provisos (Bits#(dataT, dataSz));
    VerilogEHR_1_Raw#(dataSz) ehr_raw <- mkVerilogEHRU_1_Raw;
    Reg#(dataT) ehr_ifc[1];
    
    ehr_ifc[0] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_0);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_0(pack(x));
            endmethod
        endinterface);

    return ehr_ifc;
endmodule

(* always_ready *)
interface VerilogEHR_2_Raw#(numeric type dataSz);
    method Bit#(dataSz) read_0;
    method Action write_0(Bit#(dataSz) x);
    method Bit#(dataSz) read_1;
    method Action write_1(Bit#(dataSz) x);
endinterface

import "BVI" EHR_2 =
module mkVerilogEHR_2_Raw#(Bit#(dataSz) init)(VerilogEHR_2_Raw#(dataSz));
    parameter DATA_SZ = valueOf(dataSz);
    parameter RESET_VAL = init;

    default_clock clk(CLK);
    default_reset rst(RST_N);

    method read_0 read_0;
    method write_0(write_0) enable (EN_write_0);
    method read_1 read_1;
    method write_1(write_1) enable (EN_write_1);

    // intra-port scheduling
    schedule (read_0) CF (read_0);
    schedule (read_0) SB (write_0);
    schedule (write_0) SBR (write_0);
    schedule (read_1) CF (read_1);
    schedule (read_1) SB (write_1);
    schedule (write_1) SBR (write_1);

    // inter-port scheduling
    schedule (read_0, write_0) SB (read_1, write_1);

    // paths
    path (write_0, read_1);
    path (EN_write_0, read_1);
endmodule

import "BVI" EHRU_2 =
module mkVerilogEHRU_2_Raw(VerilogEHR_2_Raw#(dataSz));
    parameter DATA_SZ = valueOf(dataSz);

    default_clock clk(CLK);
    no_reset;

    method read_0 read_0;
    method write_0(write_0) enable (EN_write_0);
    method read_1 read_1;
    method write_1(write_1) enable (EN_write_1);

    // intra-port scheduling
    schedule (read_0) CF (read_0);
    schedule (read_0) SB (write_0);
    schedule (write_0) SBR (write_0);
    schedule (read_1) CF (read_1);
    schedule (read_1) SB (write_1);
    schedule (write_1) SBR (write_1);

    // inter-port scheduling
    schedule (read_0, write_0) SB (read_1, write_1);

    // paths
    path (write_0, read_1);
    path (EN_write_0, read_1);
endmodule

module mkVerilogEHR_2#(dataT init)(VerilogEHR#(dataT)) provisos (Bits#(dataT, dataSz));
    VerilogEHR_2_Raw#(dataSz) ehr_raw <- mkVerilogEHR_2_Raw(pack(init));
    Reg#(dataT) ehr_ifc[2];
    
    ehr_ifc[0] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_0);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_0(pack(x));
            endmethod
        endinterface);
    ehr_ifc[1] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_1);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_1(pack(x));
            endmethod
        endinterface);

    return ehr_ifc;
endmodule

module mkVerilogEHRU_2(VerilogEHR#(dataT)) provisos (Bits#(dataT, dataSz));
    VerilogEHR_2_Raw#(dataSz) ehr_raw <- mkVerilogEHRU_2_Raw;
    Reg#(dataT) ehr_ifc[2];
    
    ehr_ifc[0] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_0);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_0(pack(x));
            endmethod
        endinterface);
    ehr_ifc[1] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_1);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_1(pack(x));
            endmethod
        endinterface);

    return ehr_ifc;
endmodule

(* always_ready *)
interface VerilogEHR_3_Raw#(numeric type dataSz);
    method Bit#(dataSz) read_0;
    method Action write_0(Bit#(dataSz) x);
    method Bit#(dataSz) read_1;
    method Action write_1(Bit#(dataSz) x);
    method Bit#(dataSz) read_2;
    method Action write_2(Bit#(dataSz) x);
endinterface

import "BVI" EHR_3 =
module mkVerilogEHR_3_Raw#(Bit#(dataSz) init)(VerilogEHR_3_Raw#(dataSz));
    parameter DATA_SZ = valueOf(dataSz);
    parameter RESET_VAL = init;

    default_clock clk(CLK);
    default_reset rst(RST_N);

    method read_0 read_0;
    method write_0(write_0) enable (EN_write_0);
    method read_1 read_1;
    method write_1(write_1) enable (EN_write_1);
    method read_2 read_2;
    method write_2(write_2) enable (EN_write_2);

    // intra-port scheduling
    schedule (read_0) CF (read_0);
    schedule (read_0) SB (write_0);
    schedule (write_0) SBR (write_0);
    schedule (read_1) CF (read_1);
    schedule (read_1) SB (write_1);
    schedule (write_1) SBR (write_1);
    schedule (read_2) CF (read_2);
    schedule (read_2) SB (write_2);
    schedule (write_2) SBR (write_2);

    // inter-port scheduling
    schedule (read_0, write_0) SB (read_1, write_1);
    schedule (read_0, write_0) SB (read_2, write_2);
    schedule (read_1, write_1) SB (read_2, write_2);

    // paths
    path (write_0, read_1);
    path (EN_write_0, read_1);
    path (write_0, read_2);
    path (EN_write_0, read_2);
    path (write_1, read_2);
    path (EN_write_1, read_2);
endmodule

import "BVI" EHRU_3 =
module mkVerilogEHRU_3_Raw(VerilogEHR_3_Raw#(dataSz));
    parameter DATA_SZ = valueOf(dataSz);

    default_clock clk(CLK);
    no_reset;

    method read_0 read_0;
    method write_0(write_0) enable (EN_write_0);
    method read_1 read_1;
    method write_1(write_1) enable (EN_write_1);
    method read_2 read_2;
    method write_2(write_2) enable (EN_write_2);

    // intra-port scheduling
    schedule (read_0) CF (read_0);
    schedule (read_0) SB (write_0);
    schedule (write_0) SBR (write_0);
    schedule (read_1) CF (read_1);
    schedule (read_1) SB (write_1);
    schedule (write_1) SBR (write_1);
    schedule (read_2) CF (read_2);
    schedule (read_2) SB (write_2);
    schedule (write_2) SBR (write_2);

    // inter-port scheduling
    schedule (read_0, write_0) SB (read_1, write_1);
    schedule (read_0, write_0) SB (read_2, write_2);
    schedule (read_1, write_1) SB (read_2, write_2);

    // paths
    path (write_0, read_1);
    path (EN_write_0, read_1);
    path (write_0, read_2);
    path (EN_write_0, read_2);
    path (write_1, read_2);
    path (EN_write_1, read_2);
endmodule

module mkVerilogEHR_3#(dataT init)(VerilogEHR#(dataT)) provisos (Bits#(dataT, dataSz));
    VerilogEHR_3_Raw#(dataSz) ehr_raw <- mkVerilogEHR_3_Raw(pack(init));
    Reg#(dataT) ehr_ifc[3];
    
    ehr_ifc[0] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_0);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_0(pack(x));
            endmethod
        endinterface);
    ehr_ifc[1] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_1);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_1(pack(x));
            endmethod
        endinterface);
    ehr_ifc[2] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_2);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_2(pack(x));
            endmethod
        endinterface);

    return ehr_ifc;
endmodule

module mkVerilogEHRU_3(VerilogEHR#(dataT)) provisos (Bits#(dataT, dataSz));
    VerilogEHR_3_Raw#(dataSz) ehr_raw <- mkVerilogEHRU_3_Raw;
    Reg#(dataT) ehr_ifc[3];
    
    ehr_ifc[0] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_0);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_0(pack(x));
            endmethod
        endinterface);
    ehr_ifc[1] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_1);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_1(pack(x));
            endmethod
        endinterface);
    ehr_ifc[2] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_2);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_2(pack(x));
            endmethod
        endinterface);

    return ehr_ifc;
endmodule

(* always_ready *)
interface VerilogEHR_4_Raw#(numeric type dataSz);
    method Bit#(dataSz) read_0;
    method Action write_0(Bit#(dataSz) x);
    method Bit#(dataSz) read_1;
    method Action write_1(Bit#(dataSz) x);
    method Bit#(dataSz) read_2;
    method Action write_2(Bit#(dataSz) x);
    method Bit#(dataSz) read_3;
    method Action write_3(Bit#(dataSz) x);
endinterface

import "BVI" EHR_4 =
module mkVerilogEHR_4_Raw#(Bit#(dataSz) init)(VerilogEHR_4_Raw#(dataSz));
    parameter DATA_SZ = valueOf(dataSz);
    parameter RESET_VAL = init;

    default_clock clk(CLK);
    default_reset rst(RST_N);

    method read_0 read_0;
    method write_0(write_0) enable (EN_write_0);
    method read_1 read_1;
    method write_1(write_1) enable (EN_write_1);
    method read_2 read_2;
    method write_2(write_2) enable (EN_write_2);
    method read_3 read_3;
    method write_3(write_3) enable (EN_write_3);

    // intra-port scheduling
    schedule (read_0) CF (read_0);
    schedule (read_0) SB (write_0);
    schedule (write_0) SBR (write_0);
    schedule (read_1) CF (read_1);
    schedule (read_1) SB (write_1);
    schedule (write_1) SBR (write_1);
    schedule (read_2) CF (read_2);
    schedule (read_2) SB (write_2);
    schedule (write_2) SBR (write_2);
    schedule (read_3) CF (read_3);
    schedule (read_3) SB (write_3);
    schedule (write_3) SBR (write_3);

    // inter-port scheduling
    schedule (read_0, write_0) SB (read_1, write_1);
    schedule (read_0, write_0) SB (read_2, write_2);
    schedule (read_0, write_0) SB (read_3, write_3);
    schedule (read_1, write_1) SB (read_2, write_2);
    schedule (read_1, write_1) SB (read_3, write_3);
    schedule (read_2, write_2) SB (read_3, write_3);

    // paths
    path (write_0, read_1);
    path (EN_write_0, read_1);
    path (write_0, read_2);
    path (EN_write_0, read_2);
    path (write_0, read_3);
    path (EN_write_0, read_3);
    path (write_1, read_2);
    path (EN_write_1, read_2);
    path (write_1, read_3);
    path (EN_write_1, read_3);
    path (write_2, read_3);
    path (EN_write_2, read_3);
endmodule

import "BVI" EHRU_4 =
module mkVerilogEHRU_4_Raw(VerilogEHR_4_Raw#(dataSz));
    parameter DATA_SZ = valueOf(dataSz);

    default_clock clk(CLK);
    no_reset;

    method read_0 read_0;
    method write_0(write_0) enable (EN_write_0);
    method read_1 read_1;
    method write_1(write_1) enable (EN_write_1);
    method read_2 read_2;
    method write_2(write_2) enable (EN_write_2);
    method read_3 read_3;
    method write_3(write_3) enable (EN_write_3);

    // intra-port scheduling
    schedule (read_0) CF (read_0);
    schedule (read_0) SB (write_0);
    schedule (write_0) SBR (write_0);
    schedule (read_1) CF (read_1);
    schedule (read_1) SB (write_1);
    schedule (write_1) SBR (write_1);
    schedule (read_2) CF (read_2);
    schedule (read_2) SB (write_2);
    schedule (write_2) SBR (write_2);
    schedule (read_3) CF (read_3);
    schedule (read_3) SB (write_3);
    schedule (write_3) SBR (write_3);

    // inter-port scheduling
    schedule (read_0, write_0) SB (read_1, write_1);
    schedule (read_0, write_0) SB (read_2, write_2);
    schedule (read_0, write_0) SB (read_3, write_3);
    schedule (read_1, write_1) SB (read_2, write_2);
    schedule (read_1, write_1) SB (read_3, write_3);
    schedule (read_2, write_2) SB (read_3, write_3);

    // paths
    path (write_0, read_1);
    path (EN_write_0, read_1);
    path (write_0, read_2);
    path (EN_write_0, read_2);
    path (write_0, read_3);
    path (EN_write_0, read_3);
    path (write_1, read_2);
    path (EN_write_1, read_2);
    path (write_1, read_3);
    path (EN_write_1, read_3);
    path (write_2, read_3);
    path (EN_write_2, read_3);
endmodule

module mkVerilogEHR_4#(dataT init)(VerilogEHR#(dataT)) provisos (Bits#(dataT, dataSz));
    VerilogEHR_4_Raw#(dataSz) ehr_raw <- mkVerilogEHR_4_Raw(pack(init));
    Reg#(dataT) ehr_ifc[4];
    
    ehr_ifc[0] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_0);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_0(pack(x));
            endmethod
        endinterface);
    ehr_ifc[1] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_1);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_1(pack(x));
            endmethod
        endinterface);
    ehr_ifc[2] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_2);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_2(pack(x));
            endmethod
        endinterface);
    ehr_ifc[3] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_3);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_3(pack(x));
            endmethod
        endinterface);

    return ehr_ifc;
endmodule

module mkVerilogEHRU_4(VerilogEHR#(dataT)) provisos (Bits#(dataT, dataSz));
    VerilogEHR_4_Raw#(dataSz) ehr_raw <- mkVerilogEHRU_4_Raw;
    Reg#(dataT) ehr_ifc[4];
    
    ehr_ifc[0] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_0);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_0(pack(x));
            endmethod
        endinterface);
    ehr_ifc[1] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_1);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_1(pack(x));
            endmethod
        endinterface);
    ehr_ifc[2] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_2);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_2(pack(x));
            endmethod
        endinterface);
    ehr_ifc[3] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_3);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_3(pack(x));
            endmethod
        endinterface);

    return ehr_ifc;
endmodule

(* always_ready *)
interface VerilogEHR_5_Raw#(numeric type dataSz);
    method Bit#(dataSz) read_0;
    method Action write_0(Bit#(dataSz) x);
    method Bit#(dataSz) read_1;
    method Action write_1(Bit#(dataSz) x);
    method Bit#(dataSz) read_2;
    method Action write_2(Bit#(dataSz) x);
    method Bit#(dataSz) read_3;
    method Action write_3(Bit#(dataSz) x);
    method Bit#(dataSz) read_4;
    method Action write_4(Bit#(dataSz) x);
endinterface

import "BVI" EHR_5 =
module mkVerilogEHR_5_Raw#(Bit#(dataSz) init)(VerilogEHR_5_Raw#(dataSz));
    parameter DATA_SZ = valueOf(dataSz);
    parameter RESET_VAL = init;

    default_clock clk(CLK);
    default_reset rst(RST_N);

    method read_0 read_0;
    method write_0(write_0) enable (EN_write_0);
    method read_1 read_1;
    method write_1(write_1) enable (EN_write_1);
    method read_2 read_2;
    method write_2(write_2) enable (EN_write_2);
    method read_3 read_3;
    method write_3(write_3) enable (EN_write_3);
    method read_4 read_4;
    method write_4(write_4) enable (EN_write_4);

    // intra-port scheduling
    schedule (read_0) CF (read_0);
    schedule (read_0) SB (write_0);
    schedule (write_0) SBR (write_0);
    schedule (read_1) CF (read_1);
    schedule (read_1) SB (write_1);
    schedule (write_1) SBR (write_1);
    schedule (read_2) CF (read_2);
    schedule (read_2) SB (write_2);
    schedule (write_2) SBR (write_2);
    schedule (read_3) CF (read_3);
    schedule (read_3) SB (write_3);
    schedule (write_3) SBR (write_3);
    schedule (read_4) CF (read_4);
    schedule (read_4) SB (write_4);
    schedule (write_4) SBR (write_4);

    // inter-port scheduling
    schedule (read_0, write_0) SB (read_1, write_1);
    schedule (read_0, write_0) SB (read_2, write_2);
    schedule (read_0, write_0) SB (read_3, write_3);
    schedule (read_0, write_0) SB (read_4, write_4);
    schedule (read_1, write_1) SB (read_2, write_2);
    schedule (read_1, write_1) SB (read_3, write_3);
    schedule (read_1, write_1) SB (read_4, write_4);
    schedule (read_2, write_2) SB (read_3, write_3);
    schedule (read_2, write_2) SB (read_4, write_4);
    schedule (read_3, write_3) SB (read_4, write_4);

    // paths
    path (write_0, read_1);
    path (EN_write_0, read_1);
    path (write_0, read_2);
    path (EN_write_0, read_2);
    path (write_0, read_3);
    path (EN_write_0, read_3);
    path (write_0, read_4);
    path (EN_write_0, read_4);
    path (write_1, read_2);
    path (EN_write_1, read_2);
    path (write_1, read_3);
    path (EN_write_1, read_3);
    path (write_1, read_4);
    path (EN_write_1, read_4);
    path (write_2, read_3);
    path (EN_write_2, read_3);
    path (write_2, read_4);
    path (EN_write_2, read_4);
    path (write_3, read_4);
    path (EN_write_3, read_4);
endmodule

import "BVI" EHRU_5 =
module mkVerilogEHRU_5_Raw(VerilogEHR_5_Raw#(dataSz));
    parameter DATA_SZ = valueOf(dataSz);

    default_clock clk(CLK);
    no_reset;

    method read_0 read_0;
    method write_0(write_0) enable (EN_write_0);
    method read_1 read_1;
    method write_1(write_1) enable (EN_write_1);
    method read_2 read_2;
    method write_2(write_2) enable (EN_write_2);
    method read_3 read_3;
    method write_3(write_3) enable (EN_write_3);
    method read_4 read_4;
    method write_4(write_4) enable (EN_write_4);

    // intra-port scheduling
    schedule (read_0) CF (read_0);
    schedule (read_0) SB (write_0);
    schedule (write_0) SBR (write_0);
    schedule (read_1) CF (read_1);
    schedule (read_1) SB (write_1);
    schedule (write_1) SBR (write_1);
    schedule (read_2) CF (read_2);
    schedule (read_2) SB (write_2);
    schedule (write_2) SBR (write_2);
    schedule (read_3) CF (read_3);
    schedule (read_3) SB (write_3);
    schedule (write_3) SBR (write_3);
    schedule (read_4) CF (read_4);
    schedule (read_4) SB (write_4);
    schedule (write_4) SBR (write_4);

    // inter-port scheduling
    schedule (read_0, write_0) SB (read_1, write_1);
    schedule (read_0, write_0) SB (read_2, write_2);
    schedule (read_0, write_0) SB (read_3, write_3);
    schedule (read_0, write_0) SB (read_4, write_4);
    schedule (read_1, write_1) SB (read_2, write_2);
    schedule (read_1, write_1) SB (read_3, write_3);
    schedule (read_1, write_1) SB (read_4, write_4);
    schedule (read_2, write_2) SB (read_3, write_3);
    schedule (read_2, write_2) SB (read_4, write_4);
    schedule (read_3, write_3) SB (read_4, write_4);

    // paths
    path (write_0, read_1);
    path (EN_write_0, read_1);
    path (write_0, read_2);
    path (EN_write_0, read_2);
    path (write_0, read_3);
    path (EN_write_0, read_3);
    path (write_0, read_4);
    path (EN_write_0, read_4);
    path (write_1, read_2);
    path (EN_write_1, read_2);
    path (write_1, read_3);
    path (EN_write_1, read_3);
    path (write_1, read_4);
    path (EN_write_1, read_4);
    path (write_2, read_3);
    path (EN_write_2, read_3);
    path (write_2, read_4);
    path (EN_write_2, read_4);
    path (write_3, read_4);
    path (EN_write_3, read_4);
endmodule

module mkVerilogEHR_5#(dataT init)(VerilogEHR#(dataT)) provisos (Bits#(dataT, dataSz));
    VerilogEHR_5_Raw#(dataSz) ehr_raw <- mkVerilogEHR_5_Raw(pack(init));
    Reg#(dataT) ehr_ifc[5];
    
    ehr_ifc[0] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_0);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_0(pack(x));
            endmethod
        endinterface);
    ehr_ifc[1] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_1);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_1(pack(x));
            endmethod
        endinterface);
    ehr_ifc[2] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_2);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_2(pack(x));
            endmethod
        endinterface);
    ehr_ifc[3] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_3);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_3(pack(x));
            endmethod
        endinterface);
    ehr_ifc[4] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_4);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_4(pack(x));
            endmethod
        endinterface);

    return ehr_ifc;
endmodule

module mkVerilogEHRU_5(VerilogEHR#(dataT)) provisos (Bits#(dataT, dataSz));
    VerilogEHR_5_Raw#(dataSz) ehr_raw <- mkVerilogEHRU_5_Raw;
    Reg#(dataT) ehr_ifc[5];
    
    ehr_ifc[0] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_0);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_0(pack(x));
            endmethod
        endinterface);
    ehr_ifc[1] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_1);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_1(pack(x));
            endmethod
        endinterface);
    ehr_ifc[2] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_2);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_2(pack(x));
            endmethod
        endinterface);
    ehr_ifc[3] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_3);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_3(pack(x));
            endmethod
        endinterface);
    ehr_ifc[4] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_4);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_4(pack(x));
            endmethod
        endinterface);

    return ehr_ifc;
endmodule

(* always_ready *)
interface VerilogEHR_6_Raw#(numeric type dataSz);
    method Bit#(dataSz) read_0;
    method Action write_0(Bit#(dataSz) x);
    method Bit#(dataSz) read_1;
    method Action write_1(Bit#(dataSz) x);
    method Bit#(dataSz) read_2;
    method Action write_2(Bit#(dataSz) x);
    method Bit#(dataSz) read_3;
    method Action write_3(Bit#(dataSz) x);
    method Bit#(dataSz) read_4;
    method Action write_4(Bit#(dataSz) x);
    method Bit#(dataSz) read_5;
    method Action write_5(Bit#(dataSz) x);
endinterface

import "BVI" EHR_6 =
module mkVerilogEHR_6_Raw#(Bit#(dataSz) init)(VerilogEHR_6_Raw#(dataSz));
    parameter DATA_SZ = valueOf(dataSz);
    parameter RESET_VAL = init;

    default_clock clk(CLK);
    default_reset rst(RST_N);

    method read_0 read_0;
    method write_0(write_0) enable (EN_write_0);
    method read_1 read_1;
    method write_1(write_1) enable (EN_write_1);
    method read_2 read_2;
    method write_2(write_2) enable (EN_write_2);
    method read_3 read_3;
    method write_3(write_3) enable (EN_write_3);
    method read_4 read_4;
    method write_4(write_4) enable (EN_write_4);
    method read_5 read_5;
    method write_5(write_5) enable (EN_write_5);

    // intra-port scheduling
    schedule (read_0) CF (read_0);
    schedule (read_0) SB (write_0);
    schedule (write_0) SBR (write_0);
    schedule (read_1) CF (read_1);
    schedule (read_1) SB (write_1);
    schedule (write_1) SBR (write_1);
    schedule (read_2) CF (read_2);
    schedule (read_2) SB (write_2);
    schedule (write_2) SBR (write_2);
    schedule (read_3) CF (read_3);
    schedule (read_3) SB (write_3);
    schedule (write_3) SBR (write_3);
    schedule (read_4) CF (read_4);
    schedule (read_4) SB (write_4);
    schedule (write_4) SBR (write_4);
    schedule (read_5) CF (read_5);
    schedule (read_5) SB (write_5);
    schedule (write_5) SBR (write_5);

    // inter-port scheduling
    schedule (read_0, write_0) SB (read_1, write_1);
    schedule (read_0, write_0) SB (read_2, write_2);
    schedule (read_0, write_0) SB (read_3, write_3);
    schedule (read_0, write_0) SB (read_4, write_4);
    schedule (read_0, write_0) SB (read_5, write_5);
    schedule (read_1, write_1) SB (read_2, write_2);
    schedule (read_1, write_1) SB (read_3, write_3);
    schedule (read_1, write_1) SB (read_4, write_4);
    schedule (read_1, write_1) SB (read_5, write_5);
    schedule (read_2, write_2) SB (read_3, write_3);
    schedule (read_2, write_2) SB (read_4, write_4);
    schedule (read_2, write_2) SB (read_5, write_5);
    schedule (read_3, write_3) SB (read_4, write_4);
    schedule (read_3, write_3) SB (read_5, write_5);
    schedule (read_4, write_4) SB (read_5, write_5);

    // paths
    path (write_0, read_1);
    path (EN_write_0, read_1);
    path (write_0, read_2);
    path (EN_write_0, read_2);
    path (write_0, read_3);
    path (EN_write_0, read_3);
    path (write_0, read_4);
    path (EN_write_0, read_4);
    path (write_0, read_5);
    path (EN_write_0, read_5);
    path (write_1, read_2);
    path (EN_write_1, read_2);
    path (write_1, read_3);
    path (EN_write_1, read_3);
    path (write_1, read_4);
    path (EN_write_1, read_4);
    path (write_1, read_5);
    path (EN_write_1, read_5);
    path (write_2, read_3);
    path (EN_write_2, read_3);
    path (write_2, read_4);
    path (EN_write_2, read_4);
    path (write_2, read_5);
    path (EN_write_2, read_5);
    path (write_3, read_4);
    path (EN_write_3, read_4);
    path (write_3, read_5);
    path (EN_write_3, read_5);
    path (write_4, read_5);
    path (EN_write_4, read_5);
endmodule

import "BVI" EHRU_6 =
module mkVerilogEHRU_6_Raw(VerilogEHR_6_Raw#(dataSz));
    parameter DATA_SZ = valueOf(dataSz);

    default_clock clk(CLK);
    no_reset;

    method read_0 read_0;
    method write_0(write_0) enable (EN_write_0);
    method read_1 read_1;
    method write_1(write_1) enable (EN_write_1);
    method read_2 read_2;
    method write_2(write_2) enable (EN_write_2);
    method read_3 read_3;
    method write_3(write_3) enable (EN_write_3);
    method read_4 read_4;
    method write_4(write_4) enable (EN_write_4);
    method read_5 read_5;
    method write_5(write_5) enable (EN_write_5);

    // intra-port scheduling
    schedule (read_0) CF (read_0);
    schedule (read_0) SB (write_0);
    schedule (write_0) SBR (write_0);
    schedule (read_1) CF (read_1);
    schedule (read_1) SB (write_1);
    schedule (write_1) SBR (write_1);
    schedule (read_2) CF (read_2);
    schedule (read_2) SB (write_2);
    schedule (write_2) SBR (write_2);
    schedule (read_3) CF (read_3);
    schedule (read_3) SB (write_3);
    schedule (write_3) SBR (write_3);
    schedule (read_4) CF (read_4);
    schedule (read_4) SB (write_4);
    schedule (write_4) SBR (write_4);
    schedule (read_5) CF (read_5);
    schedule (read_5) SB (write_5);
    schedule (write_5) SBR (write_5);

    // inter-port scheduling
    schedule (read_0, write_0) SB (read_1, write_1);
    schedule (read_0, write_0) SB (read_2, write_2);
    schedule (read_0, write_0) SB (read_3, write_3);
    schedule (read_0, write_0) SB (read_4, write_4);
    schedule (read_0, write_0) SB (read_5, write_5);
    schedule (read_1, write_1) SB (read_2, write_2);
    schedule (read_1, write_1) SB (read_3, write_3);
    schedule (read_1, write_1) SB (read_4, write_4);
    schedule (read_1, write_1) SB (read_5, write_5);
    schedule (read_2, write_2) SB (read_3, write_3);
    schedule (read_2, write_2) SB (read_4, write_4);
    schedule (read_2, write_2) SB (read_5, write_5);
    schedule (read_3, write_3) SB (read_4, write_4);
    schedule (read_3, write_3) SB (read_5, write_5);
    schedule (read_4, write_4) SB (read_5, write_5);

    // paths
    path (write_0, read_1);
    path (EN_write_0, read_1);
    path (write_0, read_2);
    path (EN_write_0, read_2);
    path (write_0, read_3);
    path (EN_write_0, read_3);
    path (write_0, read_4);
    path (EN_write_0, read_4);
    path (write_0, read_5);
    path (EN_write_0, read_5);
    path (write_1, read_2);
    path (EN_write_1, read_2);
    path (write_1, read_3);
    path (EN_write_1, read_3);
    path (write_1, read_4);
    path (EN_write_1, read_4);
    path (write_1, read_5);
    path (EN_write_1, read_5);
    path (write_2, read_3);
    path (EN_write_2, read_3);
    path (write_2, read_4);
    path (EN_write_2, read_4);
    path (write_2, read_5);
    path (EN_write_2, read_5);
    path (write_3, read_4);
    path (EN_write_3, read_4);
    path (write_3, read_5);
    path (EN_write_3, read_5);
    path (write_4, read_5);
    path (EN_write_4, read_5);
endmodule

module mkVerilogEHR_6#(dataT init)(VerilogEHR#(dataT)) provisos (Bits#(dataT, dataSz));
    VerilogEHR_6_Raw#(dataSz) ehr_raw <- mkVerilogEHR_6_Raw(pack(init));
    Reg#(dataT) ehr_ifc[6];
    
    ehr_ifc[0] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_0);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_0(pack(x));
            endmethod
        endinterface);
    ehr_ifc[1] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_1);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_1(pack(x));
            endmethod
        endinterface);
    ehr_ifc[2] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_2);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_2(pack(x));
            endmethod
        endinterface);
    ehr_ifc[3] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_3);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_3(pack(x));
            endmethod
        endinterface);
    ehr_ifc[4] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_4);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_4(pack(x));
            endmethod
        endinterface);
    ehr_ifc[5] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_5);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_5(pack(x));
            endmethod
        endinterface);

    return ehr_ifc;
endmodule

module mkVerilogEHRU_6(VerilogEHR#(dataT)) provisos (Bits#(dataT, dataSz));
    VerilogEHR_6_Raw#(dataSz) ehr_raw <- mkVerilogEHRU_6_Raw;
    Reg#(dataT) ehr_ifc[6];
    
    ehr_ifc[0] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_0);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_0(pack(x));
            endmethod
        endinterface);
    ehr_ifc[1] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_1);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_1(pack(x));
            endmethod
        endinterface);
    ehr_ifc[2] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_2);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_2(pack(x));
            endmethod
        endinterface);
    ehr_ifc[3] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_3);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_3(pack(x));
            endmethod
        endinterface);
    ehr_ifc[4] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_4);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_4(pack(x));
            endmethod
        endinterface);
    ehr_ifc[5] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_5);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_5(pack(x));
            endmethod
        endinterface);

    return ehr_ifc;
endmodule

(* always_ready *)
interface VerilogEHR_7_Raw#(numeric type dataSz);
    method Bit#(dataSz) read_0;
    method Action write_0(Bit#(dataSz) x);
    method Bit#(dataSz) read_1;
    method Action write_1(Bit#(dataSz) x);
    method Bit#(dataSz) read_2;
    method Action write_2(Bit#(dataSz) x);
    method Bit#(dataSz) read_3;
    method Action write_3(Bit#(dataSz) x);
    method Bit#(dataSz) read_4;
    method Action write_4(Bit#(dataSz) x);
    method Bit#(dataSz) read_5;
    method Action write_5(Bit#(dataSz) x);
    method Bit#(dataSz) read_6;
    method Action write_6(Bit#(dataSz) x);
endinterface

import "BVI" EHR_7 =
module mkVerilogEHR_7_Raw#(Bit#(dataSz) init)(VerilogEHR_7_Raw#(dataSz));
    parameter DATA_SZ = valueOf(dataSz);
    parameter RESET_VAL = init;

    default_clock clk(CLK);
    default_reset rst(RST_N);

    method read_0 read_0;
    method write_0(write_0) enable (EN_write_0);
    method read_1 read_1;
    method write_1(write_1) enable (EN_write_1);
    method read_2 read_2;
    method write_2(write_2) enable (EN_write_2);
    method read_3 read_3;
    method write_3(write_3) enable (EN_write_3);
    method read_4 read_4;
    method write_4(write_4) enable (EN_write_4);
    method read_5 read_5;
    method write_5(write_5) enable (EN_write_5);
    method read_6 read_6;
    method write_6(write_6) enable (EN_write_6);

    // intra-port scheduling
    schedule (read_0) CF (read_0);
    schedule (read_0) SB (write_0);
    schedule (write_0) SBR (write_0);
    schedule (read_1) CF (read_1);
    schedule (read_1) SB (write_1);
    schedule (write_1) SBR (write_1);
    schedule (read_2) CF (read_2);
    schedule (read_2) SB (write_2);
    schedule (write_2) SBR (write_2);
    schedule (read_3) CF (read_3);
    schedule (read_3) SB (write_3);
    schedule (write_3) SBR (write_3);
    schedule (read_4) CF (read_4);
    schedule (read_4) SB (write_4);
    schedule (write_4) SBR (write_4);
    schedule (read_5) CF (read_5);
    schedule (read_5) SB (write_5);
    schedule (write_5) SBR (write_5);
    schedule (read_6) CF (read_6);
    schedule (read_6) SB (write_6);
    schedule (write_6) SBR (write_6);

    // inter-port scheduling
    schedule (read_0, write_0) SB (read_1, write_1);
    schedule (read_0, write_0) SB (read_2, write_2);
    schedule (read_0, write_0) SB (read_3, write_3);
    schedule (read_0, write_0) SB (read_4, write_4);
    schedule (read_0, write_0) SB (read_5, write_5);
    schedule (read_0, write_0) SB (read_6, write_6);
    schedule (read_1, write_1) SB (read_2, write_2);
    schedule (read_1, write_1) SB (read_3, write_3);
    schedule (read_1, write_1) SB (read_4, write_4);
    schedule (read_1, write_1) SB (read_5, write_5);
    schedule (read_1, write_1) SB (read_6, write_6);
    schedule (read_2, write_2) SB (read_3, write_3);
    schedule (read_2, write_2) SB (read_4, write_4);
    schedule (read_2, write_2) SB (read_5, write_5);
    schedule (read_2, write_2) SB (read_6, write_6);
    schedule (read_3, write_3) SB (read_4, write_4);
    schedule (read_3, write_3) SB (read_5, write_5);
    schedule (read_3, write_3) SB (read_6, write_6);
    schedule (read_4, write_4) SB (read_5, write_5);
    schedule (read_4, write_4) SB (read_6, write_6);
    schedule (read_5, write_5) SB (read_6, write_6);

    // paths
    path (write_0, read_1);
    path (EN_write_0, read_1);
    path (write_0, read_2);
    path (EN_write_0, read_2);
    path (write_0, read_3);
    path (EN_write_0, read_3);
    path (write_0, read_4);
    path (EN_write_0, read_4);
    path (write_0, read_5);
    path (EN_write_0, read_5);
    path (write_0, read_6);
    path (EN_write_0, read_6);
    path (write_1, read_2);
    path (EN_write_1, read_2);
    path (write_1, read_3);
    path (EN_write_1, read_3);
    path (write_1, read_4);
    path (EN_write_1, read_4);
    path (write_1, read_5);
    path (EN_write_1, read_5);
    path (write_1, read_6);
    path (EN_write_1, read_6);
    path (write_2, read_3);
    path (EN_write_2, read_3);
    path (write_2, read_4);
    path (EN_write_2, read_4);
    path (write_2, read_5);
    path (EN_write_2, read_5);
    path (write_2, read_6);
    path (EN_write_2, read_6);
    path (write_3, read_4);
    path (EN_write_3, read_4);
    path (write_3, read_5);
    path (EN_write_3, read_5);
    path (write_3, read_6);
    path (EN_write_3, read_6);
    path (write_4, read_5);
    path (EN_write_4, read_5);
    path (write_4, read_6);
    path (EN_write_4, read_6);
    path (write_5, read_6);
    path (EN_write_5, read_6);
endmodule

import "BVI" EHRU_7 =
module mkVerilogEHRU_7_Raw(VerilogEHR_7_Raw#(dataSz));
    parameter DATA_SZ = valueOf(dataSz);

    default_clock clk(CLK);
    no_reset;

    method read_0 read_0;
    method write_0(write_0) enable (EN_write_0);
    method read_1 read_1;
    method write_1(write_1) enable (EN_write_1);
    method read_2 read_2;
    method write_2(write_2) enable (EN_write_2);
    method read_3 read_3;
    method write_3(write_3) enable (EN_write_3);
    method read_4 read_4;
    method write_4(write_4) enable (EN_write_4);
    method read_5 read_5;
    method write_5(write_5) enable (EN_write_5);
    method read_6 read_6;
    method write_6(write_6) enable (EN_write_6);

    // intra-port scheduling
    schedule (read_0) CF (read_0);
    schedule (read_0) SB (write_0);
    schedule (write_0) SBR (write_0);
    schedule (read_1) CF (read_1);
    schedule (read_1) SB (write_1);
    schedule (write_1) SBR (write_1);
    schedule (read_2) CF (read_2);
    schedule (read_2) SB (write_2);
    schedule (write_2) SBR (write_2);
    schedule (read_3) CF (read_3);
    schedule (read_3) SB (write_3);
    schedule (write_3) SBR (write_3);
    schedule (read_4) CF (read_4);
    schedule (read_4) SB (write_4);
    schedule (write_4) SBR (write_4);
    schedule (read_5) CF (read_5);
    schedule (read_5) SB (write_5);
    schedule (write_5) SBR (write_5);
    schedule (read_6) CF (read_6);
    schedule (read_6) SB (write_6);
    schedule (write_6) SBR (write_6);

    // inter-port scheduling
    schedule (read_0, write_0) SB (read_1, write_1);
    schedule (read_0, write_0) SB (read_2, write_2);
    schedule (read_0, write_0) SB (read_3, write_3);
    schedule (read_0, write_0) SB (read_4, write_4);
    schedule (read_0, write_0) SB (read_5, write_5);
    schedule (read_0, write_0) SB (read_6, write_6);
    schedule (read_1, write_1) SB (read_2, write_2);
    schedule (read_1, write_1) SB (read_3, write_3);
    schedule (read_1, write_1) SB (read_4, write_4);
    schedule (read_1, write_1) SB (read_5, write_5);
    schedule (read_1, write_1) SB (read_6, write_6);
    schedule (read_2, write_2) SB (read_3, write_3);
    schedule (read_2, write_2) SB (read_4, write_4);
    schedule (read_2, write_2) SB (read_5, write_5);
    schedule (read_2, write_2) SB (read_6, write_6);
    schedule (read_3, write_3) SB (read_4, write_4);
    schedule (read_3, write_3) SB (read_5, write_5);
    schedule (read_3, write_3) SB (read_6, write_6);
    schedule (read_4, write_4) SB (read_5, write_5);
    schedule (read_4, write_4) SB (read_6, write_6);
    schedule (read_5, write_5) SB (read_6, write_6);

    // paths
    path (write_0, read_1);
    path (EN_write_0, read_1);
    path (write_0, read_2);
    path (EN_write_0, read_2);
    path (write_0, read_3);
    path (EN_write_0, read_3);
    path (write_0, read_4);
    path (EN_write_0, read_4);
    path (write_0, read_5);
    path (EN_write_0, read_5);
    path (write_0, read_6);
    path (EN_write_0, read_6);
    path (write_1, read_2);
    path (EN_write_1, read_2);
    path (write_1, read_3);
    path (EN_write_1, read_3);
    path (write_1, read_4);
    path (EN_write_1, read_4);
    path (write_1, read_5);
    path (EN_write_1, read_5);
    path (write_1, read_6);
    path (EN_write_1, read_6);
    path (write_2, read_3);
    path (EN_write_2, read_3);
    path (write_2, read_4);
    path (EN_write_2, read_4);
    path (write_2, read_5);
    path (EN_write_2, read_5);
    path (write_2, read_6);
    path (EN_write_2, read_6);
    path (write_3, read_4);
    path (EN_write_3, read_4);
    path (write_3, read_5);
    path (EN_write_3, read_5);
    path (write_3, read_6);
    path (EN_write_3, read_6);
    path (write_4, read_5);
    path (EN_write_4, read_5);
    path (write_4, read_6);
    path (EN_write_4, read_6);
    path (write_5, read_6);
    path (EN_write_5, read_6);
endmodule

module mkVerilogEHR_7#(dataT init)(VerilogEHR#(dataT)) provisos (Bits#(dataT, dataSz));
    VerilogEHR_7_Raw#(dataSz) ehr_raw <- mkVerilogEHR_7_Raw(pack(init));
    Reg#(dataT) ehr_ifc[7];
    
    ehr_ifc[0] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_0);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_0(pack(x));
            endmethod
        endinterface);
    ehr_ifc[1] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_1);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_1(pack(x));
            endmethod
        endinterface);
    ehr_ifc[2] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_2);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_2(pack(x));
            endmethod
        endinterface);
    ehr_ifc[3] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_3);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_3(pack(x));
            endmethod
        endinterface);
    ehr_ifc[4] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_4);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_4(pack(x));
            endmethod
        endinterface);
    ehr_ifc[5] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_5);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_5(pack(x));
            endmethod
        endinterface);
    ehr_ifc[6] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_6);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_6(pack(x));
            endmethod
        endinterface);

    return ehr_ifc;
endmodule

module mkVerilogEHRU_7(VerilogEHR#(dataT)) provisos (Bits#(dataT, dataSz));
    VerilogEHR_7_Raw#(dataSz) ehr_raw <- mkVerilogEHRU_7_Raw;
    Reg#(dataT) ehr_ifc[7];
    
    ehr_ifc[0] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_0);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_0(pack(x));
            endmethod
        endinterface);
    ehr_ifc[1] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_1);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_1(pack(x));
            endmethod
        endinterface);
    ehr_ifc[2] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_2);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_2(pack(x));
            endmethod
        endinterface);
    ehr_ifc[3] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_3);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_3(pack(x));
            endmethod
        endinterface);
    ehr_ifc[4] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_4);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_4(pack(x));
            endmethod
        endinterface);
    ehr_ifc[5] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_5);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_5(pack(x));
            endmethod
        endinterface);
    ehr_ifc[6] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_6);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_6(pack(x));
            endmethod
        endinterface);

    return ehr_ifc;
endmodule

(* always_ready *)
interface VerilogEHR_8_Raw#(numeric type dataSz);
    method Bit#(dataSz) read_0;
    method Action write_0(Bit#(dataSz) x);
    method Bit#(dataSz) read_1;
    method Action write_1(Bit#(dataSz) x);
    method Bit#(dataSz) read_2;
    method Action write_2(Bit#(dataSz) x);
    method Bit#(dataSz) read_3;
    method Action write_3(Bit#(dataSz) x);
    method Bit#(dataSz) read_4;
    method Action write_4(Bit#(dataSz) x);
    method Bit#(dataSz) read_5;
    method Action write_5(Bit#(dataSz) x);
    method Bit#(dataSz) read_6;
    method Action write_6(Bit#(dataSz) x);
    method Bit#(dataSz) read_7;
    method Action write_7(Bit#(dataSz) x);
endinterface

import "BVI" EHR_8 =
module mkVerilogEHR_8_Raw#(Bit#(dataSz) init)(VerilogEHR_8_Raw#(dataSz));
    parameter DATA_SZ = valueOf(dataSz);
    parameter RESET_VAL = init;

    default_clock clk(CLK);
    default_reset rst(RST_N);

    method read_0 read_0;
    method write_0(write_0) enable (EN_write_0);
    method read_1 read_1;
    method write_1(write_1) enable (EN_write_1);
    method read_2 read_2;
    method write_2(write_2) enable (EN_write_2);
    method read_3 read_3;
    method write_3(write_3) enable (EN_write_3);
    method read_4 read_4;
    method write_4(write_4) enable (EN_write_4);
    method read_5 read_5;
    method write_5(write_5) enable (EN_write_5);
    method read_6 read_6;
    method write_6(write_6) enable (EN_write_6);
    method read_7 read_7;
    method write_7(write_7) enable (EN_write_7);

    // intra-port scheduling
    schedule (read_0) CF (read_0);
    schedule (read_0) SB (write_0);
    schedule (write_0) SBR (write_0);
    schedule (read_1) CF (read_1);
    schedule (read_1) SB (write_1);
    schedule (write_1) SBR (write_1);
    schedule (read_2) CF (read_2);
    schedule (read_2) SB (write_2);
    schedule (write_2) SBR (write_2);
    schedule (read_3) CF (read_3);
    schedule (read_3) SB (write_3);
    schedule (write_3) SBR (write_3);
    schedule (read_4) CF (read_4);
    schedule (read_4) SB (write_4);
    schedule (write_4) SBR (write_4);
    schedule (read_5) CF (read_5);
    schedule (read_5) SB (write_5);
    schedule (write_5) SBR (write_5);
    schedule (read_6) CF (read_6);
    schedule (read_6) SB (write_6);
    schedule (write_6) SBR (write_6);
    schedule (read_7) CF (read_7);
    schedule (read_7) SB (write_7);
    schedule (write_7) SBR (write_7);

    // inter-port scheduling
    schedule (read_0, write_0) SB (read_1, write_1);
    schedule (read_0, write_0) SB (read_2, write_2);
    schedule (read_0, write_0) SB (read_3, write_3);
    schedule (read_0, write_0) SB (read_4, write_4);
    schedule (read_0, write_0) SB (read_5, write_5);
    schedule (read_0, write_0) SB (read_6, write_6);
    schedule (read_0, write_0) SB (read_7, write_7);
    schedule (read_1, write_1) SB (read_2, write_2);
    schedule (read_1, write_1) SB (read_3, write_3);
    schedule (read_1, write_1) SB (read_4, write_4);
    schedule (read_1, write_1) SB (read_5, write_5);
    schedule (read_1, write_1) SB (read_6, write_6);
    schedule (read_1, write_1) SB (read_7, write_7);
    schedule (read_2, write_2) SB (read_3, write_3);
    schedule (read_2, write_2) SB (read_4, write_4);
    schedule (read_2, write_2) SB (read_5, write_5);
    schedule (read_2, write_2) SB (read_6, write_6);
    schedule (read_2, write_2) SB (read_7, write_7);
    schedule (read_3, write_3) SB (read_4, write_4);
    schedule (read_3, write_3) SB (read_5, write_5);
    schedule (read_3, write_3) SB (read_6, write_6);
    schedule (read_3, write_3) SB (read_7, write_7);
    schedule (read_4, write_4) SB (read_5, write_5);
    schedule (read_4, write_4) SB (read_6, write_6);
    schedule (read_4, write_4) SB (read_7, write_7);
    schedule (read_5, write_5) SB (read_6, write_6);
    schedule (read_5, write_5) SB (read_7, write_7);
    schedule (read_6, write_6) SB (read_7, write_7);

    // paths
    path (write_0, read_1);
    path (EN_write_0, read_1);
    path (write_0, read_2);
    path (EN_write_0, read_2);
    path (write_0, read_3);
    path (EN_write_0, read_3);
    path (write_0, read_4);
    path (EN_write_0, read_4);
    path (write_0, read_5);
    path (EN_write_0, read_5);
    path (write_0, read_6);
    path (EN_write_0, read_6);
    path (write_0, read_7);
    path (EN_write_0, read_7);
    path (write_1, read_2);
    path (EN_write_1, read_2);
    path (write_1, read_3);
    path (EN_write_1, read_3);
    path (write_1, read_4);
    path (EN_write_1, read_4);
    path (write_1, read_5);
    path (EN_write_1, read_5);
    path (write_1, read_6);
    path (EN_write_1, read_6);
    path (write_1, read_7);
    path (EN_write_1, read_7);
    path (write_2, read_3);
    path (EN_write_2, read_3);
    path (write_2, read_4);
    path (EN_write_2, read_4);
    path (write_2, read_5);
    path (EN_write_2, read_5);
    path (write_2, read_6);
    path (EN_write_2, read_6);
    path (write_2, read_7);
    path (EN_write_2, read_7);
    path (write_3, read_4);
    path (EN_write_3, read_4);
    path (write_3, read_5);
    path (EN_write_3, read_5);
    path (write_3, read_6);
    path (EN_write_3, read_6);
    path (write_3, read_7);
    path (EN_write_3, read_7);
    path (write_4, read_5);
    path (EN_write_4, read_5);
    path (write_4, read_6);
    path (EN_write_4, read_6);
    path (write_4, read_7);
    path (EN_write_4, read_7);
    path (write_5, read_6);
    path (EN_write_5, read_6);
    path (write_5, read_7);
    path (EN_write_5, read_7);
    path (write_6, read_7);
    path (EN_write_6, read_7);
endmodule

import "BVI" EHRU_8 =
module mkVerilogEHRU_8_Raw(VerilogEHR_8_Raw#(dataSz));
    parameter DATA_SZ = valueOf(dataSz);

    default_clock clk(CLK);
    no_reset;

    method read_0 read_0;
    method write_0(write_0) enable (EN_write_0);
    method read_1 read_1;
    method write_1(write_1) enable (EN_write_1);
    method read_2 read_2;
    method write_2(write_2) enable (EN_write_2);
    method read_3 read_3;
    method write_3(write_3) enable (EN_write_3);
    method read_4 read_4;
    method write_4(write_4) enable (EN_write_4);
    method read_5 read_5;
    method write_5(write_5) enable (EN_write_5);
    method read_6 read_6;
    method write_6(write_6) enable (EN_write_6);
    method read_7 read_7;
    method write_7(write_7) enable (EN_write_7);

    // intra-port scheduling
    schedule (read_0) CF (read_0);
    schedule (read_0) SB (write_0);
    schedule (write_0) SBR (write_0);
    schedule (read_1) CF (read_1);
    schedule (read_1) SB (write_1);
    schedule (write_1) SBR (write_1);
    schedule (read_2) CF (read_2);
    schedule (read_2) SB (write_2);
    schedule (write_2) SBR (write_2);
    schedule (read_3) CF (read_3);
    schedule (read_3) SB (write_3);
    schedule (write_3) SBR (write_3);
    schedule (read_4) CF (read_4);
    schedule (read_4) SB (write_4);
    schedule (write_4) SBR (write_4);
    schedule (read_5) CF (read_5);
    schedule (read_5) SB (write_5);
    schedule (write_5) SBR (write_5);
    schedule (read_6) CF (read_6);
    schedule (read_6) SB (write_6);
    schedule (write_6) SBR (write_6);
    schedule (read_7) CF (read_7);
    schedule (read_7) SB (write_7);
    schedule (write_7) SBR (write_7);

    // inter-port scheduling
    schedule (read_0, write_0) SB (read_1, write_1);
    schedule (read_0, write_0) SB (read_2, write_2);
    schedule (read_0, write_0) SB (read_3, write_3);
    schedule (read_0, write_0) SB (read_4, write_4);
    schedule (read_0, write_0) SB (read_5, write_5);
    schedule (read_0, write_0) SB (read_6, write_6);
    schedule (read_0, write_0) SB (read_7, write_7);
    schedule (read_1, write_1) SB (read_2, write_2);
    schedule (read_1, write_1) SB (read_3, write_3);
    schedule (read_1, write_1) SB (read_4, write_4);
    schedule (read_1, write_1) SB (read_5, write_5);
    schedule (read_1, write_1) SB (read_6, write_6);
    schedule (read_1, write_1) SB (read_7, write_7);
    schedule (read_2, write_2) SB (read_3, write_3);
    schedule (read_2, write_2) SB (read_4, write_4);
    schedule (read_2, write_2) SB (read_5, write_5);
    schedule (read_2, write_2) SB (read_6, write_6);
    schedule (read_2, write_2) SB (read_7, write_7);
    schedule (read_3, write_3) SB (read_4, write_4);
    schedule (read_3, write_3) SB (read_5, write_5);
    schedule (read_3, write_3) SB (read_6, write_6);
    schedule (read_3, write_3) SB (read_7, write_7);
    schedule (read_4, write_4) SB (read_5, write_5);
    schedule (read_4, write_4) SB (read_6, write_6);
    schedule (read_4, write_4) SB (read_7, write_7);
    schedule (read_5, write_5) SB (read_6, write_6);
    schedule (read_5, write_5) SB (read_7, write_7);
    schedule (read_6, write_6) SB (read_7, write_7);

    // paths
    path (write_0, read_1);
    path (EN_write_0, read_1);
    path (write_0, read_2);
    path (EN_write_0, read_2);
    path (write_0, read_3);
    path (EN_write_0, read_3);
    path (write_0, read_4);
    path (EN_write_0, read_4);
    path (write_0, read_5);
    path (EN_write_0, read_5);
    path (write_0, read_6);
    path (EN_write_0, read_6);
    path (write_0, read_7);
    path (EN_write_0, read_7);
    path (write_1, read_2);
    path (EN_write_1, read_2);
    path (write_1, read_3);
    path (EN_write_1, read_3);
    path (write_1, read_4);
    path (EN_write_1, read_4);
    path (write_1, read_5);
    path (EN_write_1, read_5);
    path (write_1, read_6);
    path (EN_write_1, read_6);
    path (write_1, read_7);
    path (EN_write_1, read_7);
    path (write_2, read_3);
    path (EN_write_2, read_3);
    path (write_2, read_4);
    path (EN_write_2, read_4);
    path (write_2, read_5);
    path (EN_write_2, read_5);
    path (write_2, read_6);
    path (EN_write_2, read_6);
    path (write_2, read_7);
    path (EN_write_2, read_7);
    path (write_3, read_4);
    path (EN_write_3, read_4);
    path (write_3, read_5);
    path (EN_write_3, read_5);
    path (write_3, read_6);
    path (EN_write_3, read_6);
    path (write_3, read_7);
    path (EN_write_3, read_7);
    path (write_4, read_5);
    path (EN_write_4, read_5);
    path (write_4, read_6);
    path (EN_write_4, read_6);
    path (write_4, read_7);
    path (EN_write_4, read_7);
    path (write_5, read_6);
    path (EN_write_5, read_6);
    path (write_5, read_7);
    path (EN_write_5, read_7);
    path (write_6, read_7);
    path (EN_write_6, read_7);
endmodule

module mkVerilogEHR_8#(dataT init)(VerilogEHR#(dataT)) provisos (Bits#(dataT, dataSz));
    VerilogEHR_8_Raw#(dataSz) ehr_raw <- mkVerilogEHR_8_Raw(pack(init));
    Reg#(dataT) ehr_ifc[8];
    
    ehr_ifc[0] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_0);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_0(pack(x));
            endmethod
        endinterface);
    ehr_ifc[1] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_1);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_1(pack(x));
            endmethod
        endinterface);
    ehr_ifc[2] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_2);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_2(pack(x));
            endmethod
        endinterface);
    ehr_ifc[3] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_3);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_3(pack(x));
            endmethod
        endinterface);
    ehr_ifc[4] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_4);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_4(pack(x));
            endmethod
        endinterface);
    ehr_ifc[5] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_5);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_5(pack(x));
            endmethod
        endinterface);
    ehr_ifc[6] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_6);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_6(pack(x));
            endmethod
        endinterface);
    ehr_ifc[7] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_7);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_7(pack(x));
            endmethod
        endinterface);

    return ehr_ifc;
endmodule

module mkVerilogEHRU_8(VerilogEHR#(dataT)) provisos (Bits#(dataT, dataSz));
    VerilogEHR_8_Raw#(dataSz) ehr_raw <- mkVerilogEHRU_8_Raw;
    Reg#(dataT) ehr_ifc[8];
    
    ehr_ifc[0] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_0);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_0(pack(x));
            endmethod
        endinterface);
    ehr_ifc[1] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_1);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_1(pack(x));
            endmethod
        endinterface);
    ehr_ifc[2] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_2);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_2(pack(x));
            endmethod
        endinterface);
    ehr_ifc[3] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_3);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_3(pack(x));
            endmethod
        endinterface);
    ehr_ifc[4] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_4);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_4(pack(x));
            endmethod
        endinterface);
    ehr_ifc[5] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_5);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_5(pack(x));
            endmethod
        endinterface);
    ehr_ifc[6] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_6);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_6(pack(x));
            endmethod
        endinterface);
    ehr_ifc[7] =
        (interface Reg#(dataT);
            method dataT _read;
                return unpack(ehr_raw.read_7);
            endmethod
            method Action _write(dataT x);
                ehr_raw.write_7(pack(x));
            endmethod
        endinterface);

    return ehr_ifc;
endmodule


module mkVerilogEHR#(Integer num_ports, dataT init)(VerilogEHR#(dataT)) provisos (Bits#(dataT, dataSz));
    Reg#(dataT) _ifc[num_ports];
    if (num_ports == 1) begin
        _ifc <- mkVerilogEHR_1(init);
    end else
    if (num_ports == 2) begin
        _ifc <- mkVerilogEHR_2(init);
    end else
    if (num_ports == 3) begin
        _ifc <- mkVerilogEHR_3(init);
    end else
    if (num_ports == 4) begin
        _ifc <- mkVerilogEHR_4(init);
    end else
    if (num_ports == 5) begin
        _ifc <- mkVerilogEHR_5(init);
    end else
    if (num_ports == 6) begin
        _ifc <- mkVerilogEHR_6(init);
    end else
    if (num_ports == 7) begin
        _ifc <- mkVerilogEHR_7(init);
    end else
    if (num_ports == 8) begin
        _ifc <- mkVerilogEHR_8(init);
    end else
    begin
        errorM("num_ports is too large for mkVerilogEHR");
    end
    return _ifc;
endmodule
module mkVerilogEHRU#(Integer num_ports)(VerilogEHR#(dataT)) provisos (Bits#(dataT, dataSz));
    Reg#(dataT) _ifc[num_ports];
    if (num_ports == 1) begin
        _ifc <- mkVerilogEHRU_1;
    end else
    if (num_ports == 2) begin
        _ifc <- mkVerilogEHRU_2;
    end else
    if (num_ports == 3) begin
        _ifc <- mkVerilogEHRU_3;
    end else
    if (num_ports == 4) begin
        _ifc <- mkVerilogEHRU_4;
    end else
    if (num_ports == 5) begin
        _ifc <- mkVerilogEHRU_5;
    end else
    if (num_ports == 6) begin
        _ifc <- mkVerilogEHRU_6;
    end else
    if (num_ports == 7) begin
        _ifc <- mkVerilogEHRU_7;
    end else
    if (num_ports == 8) begin
        _ifc <- mkVerilogEHRU_8;
    end else
    begin
        errorM("num_ports is too large for mkVerilogEHRU");
    end
    return _ifc;
endmodule
